module top(input clk, input [7:0] btn, output [5:0] ledc, output pwmout);

always @(posedge clk) begin
end

endmodule
