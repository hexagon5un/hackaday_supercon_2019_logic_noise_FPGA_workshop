module top(input clk, input [7:0] btn, output [5:0] led, output pwmout);

always @(posedge clk) begin
end

endmodule
